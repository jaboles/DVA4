���Z     @  +   I@      �    &                                                                                                !   �   = 	   ,          � Project@Options� -�   !�     7   |+ 	   -          � File@@Version2.1  � 1.2 =   @                                                          1   �   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Access@	 Z                   .       *       (       %       5       �       I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �0    !� BuildAll!� 0!� Read Me!�$ Copyright � 1999-2001 Jona#   ,  18 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�E H   Title , Arial ,  18 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0�    "", , , , (192,192,192), 0!�- "", ( 64, 64, 832, 832), , $   �  �� 	   -          � F1ProjectWindowsR-�   !�    �  !�  !�  !�  !�  !�  !�  !�  !�                          &     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !'   �   �� 	   -          � F1ProjectButtonsf -�   !�    �                                                          )   :   �� 	   .          � F1ProjectGlossary
 -�   !     !�  !�  !�  !�  !�  !�                                    +   bin\imagemap\!� d:\DVADev\hlp\!� _!�  !�  !�  !�  !�  !� ,    !� common!� 0!� 0!� 1!� 1!� 0!�  www.domain.com\cgi--   �   n	 	   0          � Project@OptionsHTML� -�      Read Me for DVA!� 1!�  0!�  !�  !�                       /   than Boles!�  !�  !�  !� 0!�  !�  !� 0!� 0!� No!�  !� F>   T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE FILENAME PAGE3   threats, etc. to the e-mail addresses in the DVA program gr4   oup.������Jonathan Boles��Sydney, Australia��August 2001��     ��    � 3 �� �    �    ��                   6   �)  �� 	   ,          � F1ProjectStyle2�)-�  � !�F7    Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 , 8    0 , None , !�F Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  9   20 ,  0 ,  0 ,  0 , None , !�F Normal , Arial ,  10 ,  120 :   ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�F Normal , Aria;   l ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�<   F Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,?     0 , None , !�E Title , Arial ,  18 ,  120 ,  90 ,  60 ,                                                                     WIDTH VHOBJECT0 VHOBJECT1 VHOBJECT2 VHOBJECT3              @   20 ,  0 , -1 ,  0 , None , !�E Title , Arial ,  18 ,  120 ,"     90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�E Title , Arial 2   rl����Please send questions, comments, bug reports, death Q     20 ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14 ,  1B     0 , None , !�G Heading , Arial ,  14 ,  120 ,  90 ,  60 ,C    Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,D    ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�GE    90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , ArialF   ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14 ,  120 , G    , None , !�E Title , Arial ,  18 ,  120 ,  90 ,  60 ,  20 J   �  ���-   * 1 F     � Topic@Read Me  �    �  K     �    �  ��8U     �  �� ?l     � Read Me�� N|L        �  �� 	^�     � Read Me�� 
u�     � 0 �� ��   M   9  �4 /1 /Just L /Fields /Indent 0 /Text Read Me for DVAN   �� ��  � ��/P /Just L /Fields 1�60�74��Macro �MacroArg1O    �MacroArg2 �Jump �HREF file:DVA Online.url �Anchor �TARGETP   � /Indent 0 /Text Times New Roman12��Updates and infoA   rmation are available from the website:�����1DVA Online.u`   20 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , a   , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 ,R   ding , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 S     120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub HeaT    20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 ,U    None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 , V   ing , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 ,W    120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub HeadX   20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 , Y   None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 ,  Z   ng , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , [    ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Headi\    60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14]    -1 ,  0 , None , !�G Heading , Arial ,  14 ,  120 ,  90 , ^   , !�G Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 ,_   Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None �p     20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 q   None , !�I Paragraph , Arial ,  10 ,  120 ,  90 ,  20 ,  20b   ph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , c     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�I Paragrad   ,  20 ,  0 ,  0 ,  0 , None , !�I Paragraph , Arial ,  10 ,e    0 , None , !�I Paragraph , Arial ,  10 ,  120 ,  90 ,  20 f   Heading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 , g   2 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub h    ,  20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  1i   0 , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60j   eading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  k    ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub Hl   ,  20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12m    , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 n   ading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0o   ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub Hen�    ,  0 ,  0 ,  0 , None , !�I Paragraph , Arial ,  10 ,  120�   None , !�R Bulleted List Item , Arial ,  10 ,  480 ,  90 , r   ote , Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , s    ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnt    20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnote , Arial ,  8u     0 ,  0 , None , !�G Footnote , Arial ,  8 ,  120 ,  90 , v   , !�G Footnote , Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,w    Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None x   20 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnote ,y   0 ,  0 ,  0 , None , !�O Image Paragraph , Arial ,  10 ,  1z    Image Paragraph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  {    ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�O|   0 ,  20 ,  0 ,  0 ,  0 , None , !�O Image Paragraph , Arial}    None , !�O Image Paragraph , Arial ,  10 ,  120 ,  90 ,  2~   aph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 ,    ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�O Image Paragr��    20 ,  20 ,  0 ,  0 ,  0 , None , !�R Bulleted List Item , �   Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0�     10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�E �     90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Link , Arial ,�   ,  0 , None , !�R Numbered List Item , Arial ,  10 ,  480 ,�   List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 �   480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Numbered �   ,  0 ,  0 , None , !�R Numbered List Item , Arial ,  10 ,  �   ered List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 �   0 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Numb�   ,  0 ,  0 ,  0 , None , !�R Numbered List Item , Arial ,  1�    Bulleted List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 �    ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R�     20 ,  0 ,  0 ,  0 , None , !�R Bulleted List Item , Arial�   , !�R Bulleted List Item , Arial ,  10 ,  480 ,  90 ,  20 ,�   Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None �    , None , !�E Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,�    ,  20 ,  0 ,  0 ,  0 , None , !�E Index , Arial ,  10 ,  1�    0 ,  0 , None , !�E Index , Arial ,  10 ,  120 ,  90 ,  20�    , !�E Index , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �    Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None�     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Index ,�   20 ,  20 ,  10 ,  0 ,  0 , None , !�E Index , Arial ,  10 ,�   ,  0 , None , !�K Image Link , Arial ,  10 ,  120 ,  90 ,  �   age Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 �   10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�K Im�   0 ,  20 ,  10 ,  0 ,  0 , None , !�K Image Link , Arial ,  �     0 , None , !�K Image Link , Arial ,  10 ,  120 ,  90 ,  2�   ge Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,�   0 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�K Ima�    ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�E Link , Arial ,  1�     10 ,  0 ,  0 , None , !�E Link , Arial ,  10 ,  120 ,  90�   20 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�M Index Head�   l ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !��     20 ,  0 , -1 ,  0 , None , !�S Glossary Definition , Aria�   None , !�M Glossary Term , Arial ,  12 ,  120 ,  90 ,  20 ,�   rm , Arial ,  12 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , �   0 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Glossary Te�    0 , -1 ,  0 , None , !�M Glossary Term , Arial ,  12 ,  12�   !�M Glossary Term , Arial ,  12 ,  120 ,  90 ,  20 ,  20 , �   ial ,  12 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , �    ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Glossary Term , Ar�    ,  0 , None , !�M Index Heading , Arial ,  14 ,  120 ,  90�   ex Heading , Arial ,  14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1�   14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Ind�   ,  20 ,  0 , -1 ,  0 , None , !�M Index Heading , Arial ,  �    None , !�M Index Heading , Arial ,  14 ,  120 ,  90 ,  20 �   ing , Arial ,  14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 ,B�   S Glossary Definition , Arial ,  10 ,  120 ,  90 ,  20 ,  2�   ,  120 ,  90 ,  20 ,  20 ,  5 ,  0 ,  0 , None , !�P Button�   ,  5 ,  0 ,  0 , None , !�P Button Bar , Courier New ,  10 �   �P Button Bar , Courier New ,  10 ,  120 ,  90 ,  20 ,  20 �   al ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�   60 ,  20 ,  0 , -1 ,  0 , None , !�P Glossary Heading , Ari�    None , !�P Glossary Heading , Arial ,  14 ,  120 ,  90 ,  �   ing , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 ,�   ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�P Glossary Head�   -1 ,  0 , None , !�P Glossary Heading , Arial ,  14 ,  120 �   sary Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , �   0 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�P Glos�     0 ,  0 ,  0 , None , !�S Glossary Definition , Arial ,  1�   lossary Definition , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,�     10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�S G�   0 ,  0 ,  0 ,  0 , None , !�S Glossary Definition , Arial ,F�    Bar , Courier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  5 ,  0�   ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline Node �   0 ,  0 ,  0 , None , !�L Outline Node , Arial ,  10 ,  120 �   !�L Outline Node , Arial ,  10 ,  120 ,  90 ,  10 ,  10 ,  �   ial ,  10 ,  120 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , �   0 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline Node , Ar�    0 ,  0 , None , !�L Outline Node , Arial ,  10 ,  120 ,  9�    , !�E Table , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �    Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None�     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Table ,�    20 ,  20 ,  0 ,  0 ,  0 , None , !�E Table , Arial ,  10 ,�    ,  0 ,  0 , None , !�E Table , Arial ,  10 ,  120 ,  90 , �   one , !�E Table , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0�   urier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  5 ,  0 ,  0 , N�    90 ,  20 ,  20 ,  5 ,  0 ,  0 , None , !�P Button Bar , Co�    ,  0 , None , !�P Button Bar , Courier New ,  10 ,  120 , ��   , Arial ,  10 ,  120 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , Non�   , None , !�C Image , Arial ,  10 ,  120 ,  90 ,  0 ,  0 ,  �    Image , Arial ,  10 ,  120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 �    ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�C�    ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�D Line , Arial�   ,  20 ,  0 ,  0 ,  0 , None , !�D Line , Arial ,  10 ,  120�    0 ,  0 , None , !�D Line , Arial ,  10 ,  120 ,  90 ,  20 �   e , !�D Line , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �   , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , Non�    ,  440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�D Line �     10 ,  0 ,  0 ,  0 , None , !�L Outline Leaf , Arial ,  10�    None , !�L Outline Leaf , Arial ,  10 ,  440 ,  90 ,  10 ,�   eaf , Arial ,  10 ,  440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 ,�   440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline L�    ,  0 ,  0 ,  0 , None , !�L Outline Leaf , Arial ,  10 ,  �   e , !�L Outline Leaf , Arial ,  10 ,  440 ,  90 ,  10 ,  10�   0 ,  0 ,  0 , None , !�C Image , Arial ,  10 ,  120 ,  90 ,�    20 ,  20 ,  0 ,  0 ,  0 , None , !�Q Mono Spaced , Courier�    None , !�Q Mono Spaced , Courier New ,  10 ,  120 ,  90 , �   Courier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 ,�     90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�Q Mono Spaced , �    ,  0 , None , !�Q Mono Spaced , Courier New ,  10 ,  120 ,�   ect , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0�    120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Form Obj�    ,  0 ,  0 , None , !�R Form Object , MS Sans Serif ,  8 , �   m Object , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20 ,  0�    8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R For�    ,  0 ,  0 ,  0 , None , !�R Form Object , MS Sans Serif , �   R Form Object , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20�   ial ,  10 ,  120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��    120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�C Image , Ar�     0 ,  0 ,  0 ,  0 ,  0 , None , !�C Image , Arial ,  10 ,     New ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None ,                                                               �                                                              �                                                              �                                                              �                                                              �                                                                   !�  !� T�0�Read Me�Read Me� �                           �   W   �� 	   1          � F1ProjectContentList$ -�      �  !�  !�  !�  !�  !�  !�  !�  !�                          �   Index", ( 511, 0, 511, 1023), , , (192,192,192), 0!�  !�  !�   4 "Glossary", ( 0, 0, 511, 1023), , , (192,192,192), 0!�3 "�   192), 0!�. "", ( 0, 511, 1023, 511), , , (192,192,192), 0!��   , (192,192,192), 0!�, "", ( 0, 0, 1023, 511), , , (192,192,    20 ,  0 ,  0 ,  0 , None , !�                              �    !�Q Mono Spaced , Courier New ,  10 ,  120 ,  90 ,  20 ,  