���Z     @  f   I�      q   &                                       �'    �                                                     !   �   �h 	   ,          � Project@Options� -�   !�     7   |+ 	   -          � File@@Version2.1  � 1.2 �   �                                                          �   �  TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule Access ' �                  .       *       (       %       #             +      !l      %N      1V      2      <p      =�      A�      E�      gl      l�      t�      ��      ��      ��      �.      ��      ��      ��      �q      �w      �%      �'      �      ��      �C      �X      �m      ��      �F      �      ŀ      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      n0    !� BuildAll!� 0!�	 About DVA!�$ Copyright � 1999-2001 Jo1    Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 , "   �)  �� 	   ,          � F1ProjectStyle2�)-�  � !�F    "", , , , (192,192,192), 0!�- "", ( 64, 64, 832, 832), , $   �  �t 	   -          � F1ProjectWindows�-�   !�    �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�                  &     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !'   �   - 	   -          � F1ProjectButtonsn -�   !�    �                                                          )   :   �� 	   .          � F1ProjectGlossary
 -�   !     !�  !�  !�  !�  !�  !�                                    +   bin\imagemap\!� d:\DVADev\hlp\!� _!�  !�  !�  !�  !�  !� ,    !� common!� 0!� 0!� 1!� 1!� 0!�  www.domain.com\cgi--   �   n	 	   0          � Project@OptionsHTML� -�       DVA Help!� 1!�  0!�  !�  !�                            /   nathan Boles!�  !�  !�  !� 0!�  !�  !� 0!� 0!� No!�  !�@    0 , None , !�F Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  A     0 , None , !�G Heading , Arial ,  14 ,  120 ,  90 ,  60 ,2    Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,3    ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G4    90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , Arial5   ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14 ,  120 , 6    , None , !�E Title , Arial ,  18 ,  120 ,  90 ,  60 ,  20 7   Title , Arial ,  18 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  08   ,  18 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�E 9     90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�E Title , Arial :   20 ,  0 , -1 ,  0 , None , !�E Title , Arial ,  18 ,  120 ,;     0 , None , !�E Title , Arial ,  18 ,  120 ,  90 ,  60 ,  <   F Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,=   l ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�>   ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�F Normal , Aria?   20 ,  0 ,  0 ,  0 , None , !�F Normal , Arial ,  10 ,  120 nP     20 ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14 ,  1Q   ding , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 B     120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub HeaC    20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 ,D    None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 , E   ing , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 ,F    120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub HeadG   20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 , H   None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 ,  I   ng , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , J    ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G HeadiK    60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14L    -1 ,  0 , None , !�G Heading , Arial ,  14 ,  120 ,  90 , M   , !�G Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 ,N   Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None O   20 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , `   , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 ,a   ph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , R     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�I ParagraS   ,  20 ,  0 ,  0 ,  0 , None , !�I Paragraph , Arial ,  10 ,T    0 , None , !�I Paragraph , Arial ,  10 ,  120 ,  90 ,  20 U   Heading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 , V   2 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub W    ,  20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  1X   0 , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60Y   eading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  Z    ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub H[   ,  20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12\    , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 ]   ading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0^   ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub He_     20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 np   None , !�I Paragraph , Arial ,  10 ,  120 ,  90 ,  20 ,  20q   ote , Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , b    ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnc    20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnote , Arial ,  8d     0 ,  0 , None , !�G Footnote , Arial ,  8 ,  120 ,  90 , e   , !�G Footnote , Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,f    Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None g   20 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnote ,h   0 ,  0 ,  0 , None , !�O Image Paragraph , Arial ,  10 ,  1i    Image Paragraph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  j    ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�Ok   0 ,  20 ,  0 ,  0 ,  0 , None , !�O Image Paragraph , Ariall    None , !�O Image Paragraph , Arial ,  10 ,  120 ,  90 ,  2m   aph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 ,n    ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�O Image Paragro    ,  0 ,  0 ,  0 , None , !�I Paragraph , Arial ,  10 ,  1202�   None , !�R Bulleted List Item , Arial ,  10 ,  480 ,  90 , �     10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�E r     90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Link , Arial ,s   ,  0 , None , !�R Numbered List Item , Arial ,  10 ,  480 ,t   List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 u   480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Numbered v   ,  0 ,  0 , None , !�R Numbered List Item , Arial ,  10 ,  w   ered List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 x   0 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Numby   ,  0 ,  0 ,  0 , None , !�R Numbered List Item , Arial ,  1z    Bulleted List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 {    ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R|     20 ,  0 ,  0 ,  0 , None , !�R Bulleted List Item , Arial}   , !�R Bulleted List Item , Arial ,  10 ,  480 ,  90 ,  20 ,~   Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None     20 ,  20 ,  0 ,  0 ,  0 , None , !�R Bulleted List Item , ��   Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0�    0 ,  0 , None , !�E Index , Arial ,  10 ,  120 ,  90 ,  20�    , !�E Index , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �    Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None�     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Index ,�   20 ,  20 ,  10 ,  0 ,  0 , None , !�E Index , Arial ,  10 ,�   ,  0 , None , !�K Image Link , Arial ,  10 ,  120 ,  90 ,  �   age Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 �   10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�K Im�   0 ,  20 ,  10 ,  0 ,  0 , None , !�K Image Link , Arial ,  �     0 , None , !�K Image Link , Arial ,  10 ,  120 ,  90 ,  2�   ge Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,�   0 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�K Ima�    ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�E Link , Arial ,  1�     10 ,  0 ,  0 , None , !�E Link , Arial ,  10 ,  120 ,  90�    , None , !�E Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,�    ,  20 ,  0 ,  0 ,  0 , None , !�E Index , Arial ,  10 ,  1�     20 ,  0 , -1 ,  0 , None , !�S Glossary Definition , Aria�   None , !�M Glossary Term , Arial ,  12 ,  120 ,  90 ,  20 ,�   rm , Arial ,  12 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , �   0 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Glossary Te�    0 , -1 ,  0 , None , !�M Glossary Term , Arial ,  12 ,  12�   !�M Glossary Term , Arial ,  12 ,  120 ,  90 ,  20 ,  20 , �   ial ,  12 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , �    ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Glossary Term , Ar�    ,  0 , None , !�M Index Heading , Arial ,  14 ,  120 ,  90�   ex Heading , Arial ,  14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1�   14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Ind�   ,  20 ,  0 , -1 ,  0 , None , !�M Index Heading , Arial ,  �    None , !�M Index Heading , Arial ,  14 ,  120 ,  90 ,  20 �   ing , Arial ,  14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 ,�   20 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�M Index Head��   l ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !��   ,  5 ,  0 ,  0 , None , !�P Button Bar , Courier New ,  10 �   �P Button Bar , Courier New ,  10 ,  120 ,  90 ,  20 ,  20 �   al ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�   60 ,  20 ,  0 , -1 ,  0 , None , !�P Glossary Heading , Ari�    None , !�P Glossary Heading , Arial ,  14 ,  120 ,  90 ,  �   ing , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 ,�   ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�P Glossary Head�   -1 ,  0 , None , !�P Glossary Heading , Arial ,  14 ,  120 �   sary Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , �   0 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�P Glos�     0 ,  0 ,  0 , None , !�S Glossary Definition , Arial ,  1�   lossary Definition , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,�     10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�S G�   0 ,  0 ,  0 ,  0 , None , !�S Glossary Definition , Arial ,�   S Glossary Definition , Arial ,  10 ,  120 ,  90 ,  20 ,  2�   ,  120 ,  90 ,  20 ,  20 ,  5 ,  0 ,  0 , None , !�P Button�   0 ,  0 ,  0 , None , !�L Outline Node , Arial ,  10 ,  120 �   !�L Outline Node , Arial ,  10 ,  120 ,  90 ,  10 ,  10 ,  �   ial ,  10 ,  120 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , �   0 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline Node , Ar�    0 ,  0 , None , !�L Outline Node , Arial ,  10 ,  120 ,  9�    , !�E Table , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �    Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None�     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Table ,�    20 ,  20 ,  0 ,  0 ,  0 , None , !�E Table , Arial ,  10 ,�    ,  0 ,  0 , None , !�E Table , Arial ,  10 ,  120 ,  90 , �   one , !�E Table , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0�   urier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  5 ,  0 ,  0 , N�    90 ,  20 ,  20 ,  5 ,  0 ,  0 , None , !�P Button Bar , Co�    ,  0 , None , !�P Button Bar , Courier New ,  10 ,  120 , �    Bar , Courier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  5 ,  0n�   ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline Node �    Image , Arial ,  10 ,  120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 �    ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�C�    ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�D Line , Arial�   ,  20 ,  0 ,  0 ,  0 , None , !�D Line , Arial ,  10 ,  120�    0 ,  0 , None , !�D Line , Arial ,  10 ,  120 ,  90 ,  20 �   e , !�D Line , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �   , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , Non�    ,  440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�D Line �     10 ,  0 ,  0 ,  0 , None , !�L Outline Leaf , Arial ,  10�    None , !�L Outline Leaf , Arial ,  10 ,  440 ,  90 ,  10 ,�   eaf , Arial ,  10 ,  440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 ,�   440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline L�    ,  0 ,  0 ,  0 , None , !�L Outline Leaf , Arial ,  10 ,  �   e , !�L Outline Leaf , Arial ,  10 ,  440 ,  90 ,  10 ,  10�   , Arial ,  10 ,  120 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , Non�   , None , !�C Image , Arial ,  10 ,  120 ,  90 ,  0 ,  0 ,  �    None , !�Q Mono Spaced , Courier New ,  10 ,  120 ,  90 , �   Courier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 ,�     90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�Q Mono Spaced , �    ,  0 , None , !�Q Mono Spaced , Courier New ,  10 ,  120 ,�   ect , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0�    120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Form Obj�    ,  0 ,  0 , None , !�R Form Object , MS Sans Serif ,  8 , �   m Object , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20 ,  0�    8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R For�    ,  0 ,  0 ,  0 , None , !�R Form Object , MS Sans Serif , �   R Form Object , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20�   ial ,  10 ,  120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��    120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�C Image , Ar�     0 ,  0 ,  0 ,  0 ,  0 , None , !�C Image , Arial ,  10 , �   0 ,  0 ,  0 , None , !�C Image , Arial ,  10 ,  120 ,  90 ,n�    20 ,  20 ,  0 ,  0 ,  0 , None , !�Q Mono Spaced , Courier�   4 "Glossary", ( 0, 0, 511, 1023), , , (192,192,192), 0!�3 "�   Index", ( 511, 0, 511, 1023), , , (192,192,192), 0!�  !�  !�  �  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  �   ation see the DVA program group.��ICQ: 140329012����All �   Boles 1999-2001. ��All rights reserved.��For contact informT                                                               WIDTH VHOBJECT0 VHOBJECT1 VHOBJECT2 VHOBJECT3 VHOBJECT4 VHO�   omputer program is protected by copyright law. Unauthorised�   e at: 2www.railpage.org.au/railwavs. ����Warning: This c�   T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE FILENAME PAGE�   l, Paul McCabe and Winston Yang.��Visit the Railwavs websit�   sounds included with DVA are copyright Glenn Jackson-Bethel    20 ,  0 ,  0 ,  0 , None , !�                              �    !�Q Mono Spaced , Courier New ,  10 ,  120 ,  90 ,  20 ,  �    New ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None ,��   192), 0!�. "", ( 0, 511, 1023, 511), , , (192,192,192), 0!��   ut DVA�� 

;    � 0 ��y  3  �. /1 /Just L /Fields /�   Indent 0 /Text About DVA��3�  ^ �Y/P /Just L /Field�   s 1�156�163��Macro �MacroArg1 �MacroArg2 �Jump �HREF http:��   �www.icq.com �Anchor �TARGET�2�293�320��Macro �MacroArg1 �M�   acroArg2 �Jump �HREF http:��www.railpage.org.au�railwavs �A�   nchor �TARGET� /Indent 0 /Text Times New Roman12��DVA�   ��Digital Voice Announcer ��Version 4 ��Copyright Jonathan   , and will be prosecuted to the maximum extent possible und�   on of it, may result in severe civil and criminal penalties�    reproduction or distribution of this program, or any porti�   ields /Indent 0 /Text Times New Roman12��DVA stands f�   or Digital Voice Announcement. It is a program which lets y�   ou create announcements as used at CityRail stations all ov  er Sydney. The DVA distribution package consists of the act�   , (192,192,192), 0!�, "", ( 0, 0, 1023, 511), , , (192,192,*�   �� A    �	 About DVA�� �    �  �� 	�*    �	 Abo,   DVA�� �!� T�1�What is DVA?�What is DVA� �!�( T�1�Past Dev   !�  !� T�0�About DVA�About DVA� �!� F�0�Introduction to  H  � 	   1          � F1ProjectContentList-�      er the law. ����D�    � 3 ���    �   ��      ����- <  . 5 J     � Topic@What is DVA  �       �    �                                             ds) in places such as shopping centres or theatres. ����   any public address system (provided you have the right soun	  urce files to get you started. DVA can also be used to run 
  ual DVA program, hundreds of CityRail sounds, and sample so   �    �    �  ��<Y     �  �� Cu     � What is DV  A?�� R�     �  �� 	b�     � Printing a File�� 
~�       � 0 �� ��     � 3 �� �  6  �1 /1 /Just L /Fields �   /Indent 0 /Text What is DVA?�� ��  � ��/P /Just L /F  /LMargin /TMargin /RMargin /BMargin /Meta ��:�     �  "  ckImage /Fixed /Sound /Loop /Base /Isindex /Prompt /Center !  ust L /Fields /Indent 0 /Text Times New Roman12��The   st L /Stack Y /Indent 0 /Width /Height�� �(  �  �� /P /J  �     � 0 �� ��   8  �3 /1 /Just L /Fields /Indent 0 /Te  xt Opening a File�� ��  �  �� /P /Just L /Fields /Inde  nt 0 /Text Times New Roman12��Opening a file places i  t in the editing area. From there you can edit, play, or co  mpile it. DVA can open MVA files as well as DVA Files.����   �  ?  �: /4 /Just L /Fields /Indent 0 /Text 11To Ope  n a File:���� �  o  �j /B /Just L /Fields /Indent 0 /T  ext In Windows Explorer, simply right-click the file and thE  BJECT5 VHOBJECT6 VHOBJECT7 VHOBJECT8 VHOBJECT9 VHOBJECT10 V  en click Open.����  E  �@ /P /Just L /Fields /Indent 8  0 /Text Times New Roman12��OR��%%  4  �/ /E /Ju     ���- �  , 3 �     � Topic@About DVA  �    �      �  �  �� /Color1 /Color2 /Color3 /Color4 /Color5 /Ba0  Options menu (shortcut Alt+O) contains commands for cha1  come a long way from its roots. Development began in 1999 w"  .quickbasic.net �Anchor �TARGET� /Indent 0 /Text ��DVA has #  �228��Macro �MacroArg1 �MacroArg2 �Jump �HREF http:��qb4all$  F http:��www.basicguru.com�abc�rapidq �Anchor �TARGET�2�219%  L /Fields 1�346�352��Macro �MacroArg1 �MacroArg2 �Jump �HRE&  /Indent 0 /Text Past Development�� �D  . �)/P /Just '    � 0 �� ��     � 3 �� �  :  �5 /1 /Just L /Fields (  Development�� W�     �  �� 	g�     � Topic1�� 
��   )      �    �    �  ��A^     �  �� H~     � Past *  ]  j��- !  3 : O     � Topic@Past Development  �\  elopment�Past Development� �!�  T�1�New in DVA 4�New in DVA      � 5 ��1�    �   ��                           -  ialog box for changing many of DVA's settings.���� ��  .  /Indent 0 /Text Preferences... displays the Preferences d/  nging DVA's settings: ���� ��  �  �~ /B /Just L /Fields @  ith the concept of DVA being realised in the form of an MS-A   can open a file by double-clicking it.����    � 10 �2   If you have specified so in Options, Preferences, you3  ����.�  �  �� /P /Just L /Fields /Indent 0 /Text Note:4   /Text Browse for the file, select it, and then click OK.5  ess Ctrl+O.������  ^  �Y /E /Just L /Fields /Indent 06   /Just L /Fields /Indent 0 /Text Click File, Open or pr7  st L /Fields /Indent 0 /Text Start DVA.������  Q  �L /E    y been a 'great leap forward'. ���� �T    �    M9  ed and advanced version to date; each new version has reall:  ew features added and hence this version is the most enhanc;  d has reached version number 4. Each new version has seen n<  major version numbers. Now DVA is written in 1Rapid-Q an=  l, and Turbo Pascal for Windows and has been through three >  ough the hands of MS-DOS Batch, 2QuickBasic, Turbo Pasca?  DOS batch file. Since then, until today, DVA has passed thr    ��    �   ��                                   C  Create a New File:���� �;  �  �� /B /Just L /Fields /InD  dent 0 /Text From a Windows Explorer window, simply right-cF  lick in a blank area, point to New, then click DVA SourcU  HOBJECT11 VHOBJECT12 VHOBJECT13 VHOBJECT14 VHOBJECT15 VHOBJG  e. Then you can open the file for editing.�� �  E  �@ H  /P /Just L /Fields /Indent 0 /Text Times New Roman12��I  OR��}�  4  �/ /E /Just L /Fields /Indent 0 /Text StaJ  rt DVA.����D$  O  �J /E /Just L /Fields /Indent 0 /TextK   Click File, New, or press Ctrl+N.���5    � 7 �    ��E    �   ->                                   �  ndent 0 /Text Printing a File�� ��  �  �� /P /Just L /�  le� �!�" T�1�Saving a File�Saving a File� �!�& T�1�PrintingO  �  ]w��B 1  1 8 M     � Topic@Opening a File  �  P    �    �    �  ��?\     �  �� Fz     � Opening   a File�� U�     �  �� 	e�     � Opening a File�� 
�nB  Just L /Fields /Indent 0 /Text Times New Roman��11To S  tion point. �����$  ^  �Y /B /Just L /Fields /Indent 0 W  /Text Clear (shortcut Del) deletes the selected text. �                                                               y  ECT16 VHOBJECT17 VHOBJECT18 VHOBJECT19 VHOBJECT20 VHOBJECT2]  N  ���9 2  6 = R     � Topic@Creating a New FileX  ���9�  q  �l /B /Just L /Fields /Indent 0 /Text Select�   All (shortcut Ctrl+A) Selects all text in the editing aZ  tions Menu�� ��  �  �� /I /Jump /Link j:\HLP\WINHELP4\S  OURCE\COMMON\OPTION~1.BMP /Macro /Play /Popup /Border 0 /JuM  e�Creating a New File� �!�$ T�1�Opening a File�Opening a Fi[   4� �!� F�0�Tasks/Procedures�� �!�. T�1�Creating a New Fil^    �    �    �    �  ��Da     �  �� K�     � Cr_  eating a New File�� Z�     �  �� 	j�     � Creating a`   New File�� 
��     � 0 �� �  =  �8 /1 /Just L /FieldQ  s /Indent 0 /Text Creating a New File�� �t  Y  �T /4 /�R  ut Ctrl+V) Inserts any text in the clipboard at the inserq  DOS program to play its sounds. The newer way to play is mub  sound files. In previous versions, it launched an external c  L /Fields /Indent 0 /Text DVA now uses Windows to play its d  dent 0 /Text ��Enhanced Playback�� 	  ? �:/P /Just e  rsion. Here they are:�� ȼ  =  �8 /4 /Just L /Fields /Inf  Indent 0 /Text ��DVA has many new features in its latest veg   0 /Text New in DVA 4�� �t  i  �d /P /Just L /Fields /h  �� ��     � 19 �� �   6  �1 /1 /Just L /Fields /Indenti  A 4�� S�     �  �� 	c�     � Topic1�� 
�     � 0 j    �    �    �  ��=Z     �  �� Dv     � New in DVk  ;  �+��] %  / 6 K     � Topic@New in DVA 4  �  L   � 0 �� ��     � 5 �� �  9  �4 /1 /Just L /Fields /Im  ng a File�� V�     �  �� 	f�     � Topic1�� 
��    n     �    �    �  ��@]     �  �� G|     � Printio    4���3 =  2 9 N     � Topic@Printing a File  � n�  ch faster and more bug-free, since it is built right into W�  t As well as writing your files in the the normal way with r   List Box����   �/P /Just L /Fields /Indent 0 /Texs  D�  >  �9 /4 /Just L /Fields /Indent 0 /Text Quick-Buildt  nding a string of text, and searching-and-replacing. ����u   the DVA program. The DVA program now has facilities for fiv  .00, you can now edit DVA (and MVA) files right from withinw    �  �� /P /Just L /Fields /Indent 0 /Text As of version 4x  /Indent 0 /Text Full-featured Built-in Text Editor��c�y  s in too low quality. �����  L  �G /4 /Just L /Fields z  a slow computer and playing the file through Windows result{   an MS-DOS batch file. You may want to do this if you have |   L /Fields /Indent 0 /Text DVA now allows you to compile to}  t Compile to an MS-DOS Batch File���;  �  �� /P /Just~   now... ����}Z  I  �D /4 /Just L /Fields /Indent 0 /Tex  indows. Of course, if you want to play the old way, you can��  the built in editor, you can very quickly create your files�  ening, playing, or compiling a file, and you can specify wh�   also customisable. There are right-click menu items for op�  lds /Indent 0 /Text DVA includes shell integration which is�  ble 100% Shell Integration ��-(
   �/P /Just L /Fie�  ��	  N  �I /4 /Just L /Fields /Indent 0 /Text Customisa�  n DVA. DVA lets you open, save and print any MVA file. ����  ndent 0 /Text You can now play and compile your MVA files i�  /Text MVA-Compatible��ӽ  �  �� /P /Just L /Fields /I�  e are used. �����$  8  �3 /4 /Just L /Fields /Indent 0 �  est the file, since only files that are there and accessibl�   create a DVA or MVA file. It also eliminates the need to t�  t the insertion point. This makes it very quick and easy to�   Simply double click a file to add it to the editing area a�  s box contains every file in your default sounds directory.�   with the list box appearing at the side of the window. Thi*�  ich action is the default, for when the file is double-clic�    �    �    �  ��>[     �  �� Ex     � Saving a    d.��
�2    �   � +                               �  ity now means that this requirement is completely eliminate�   all the sounds to play correctly. DVA's Windows compatibil�  filename support meant that an index file was mandatory for�  need for an index file. In previous versions, lack of long �   L /Fields /Indent 0 /Text Version 4 of DVA eliminates the �  ent 0 /Text Index File Eliminated��
{"  6 �1/P /Just�   are implemented. ����	1�  ?  �: /4 /Just L /Fields /Ind�  onsistent dialogs for operations such as opening and saving�  hare text on the clipboard, use long filenames, and fully c�  it compiler, it is compatible fully with Windows. You can s�  ndent 0 /Text Because DVA is now written in Rapid-Q, a 32-b�  Windows Compatibility���   �/P /Just L /Fields /I�  ked. �����r
  ?  �: /4 /Just L /Fields /Indent 0 /Text n�   File�� T�     �  �� 	d�     � Saving a File�� 
��  �  the text box����49  8  �3 /E /Just L /Fields /Indent 0 �  t Choose the format (.dva or .mva) and enter a new name in �  As.... ������  o  �j /E /Just L /Fields /Indent 0 /Tex�   �A /E /Just L /Fields /Indent 0 /Text Click File, Save �  le with a new name or in a different format:����c|  F �   h  �c /4 /Just L /Fields /Indent 0 /Text 11To save a fi�   /Text Press Ctrl+S, or click File, Save. �����+ �  usly saved: ���� �  S  �N /B /Just L /Fields /Indent 0�  s /Indent 0 /Text 11To save a file which you have previo�   Save As... dialog box. ���� �Z  `  �[ /4 /Just L /Field�  ed.dva. Any save command will automatically take you to the�  ile and have not saved it yet, it will have the name Untitl�   /Text Times New Roman12��If you have created a new f�  Saving a File�� ��  �  �� /P /Just L /Fields /Indent 0�     � 0 �� ��   7  �2 /1 /Just L /Fields /Indent 0 /Text ��  /Text Click Save. �����J    � 9 ���Z    �   �    �    �    �  ��?\     �  �� Fz     � Playing�  �  W���? A  1 8 M     � Topic@Playing a File  �  �   a File�Printing a File� �!�$ T�1�Playing a File�Playing a L  File� �!�( T�1�Compiling a File�Compiling a File� �!� F�0�    ftware.org �����h    �   ba                       '.���    �   .                               �   in Options, Preferences. The default setting is 'LPT1:�   DVA source will be printed to the device or file specified�  dent 0 /Text Press Ctrl+P, or click File, Print. Your�  To Print a File:���� �  �  �� /B /Just L /Fields /In�  . ���� �%  A  �< /4 /Just L /Fields /Indent 0 /Text 11�  m. You can set this device/file in Options, Preferences�   network printer/device, and also to any file on your syste�  Fields /Indent 0 /Text ��DVA lets you print to any local or    BS                                                     *�   a File�� U�     �  �� 	e�     � Topic1�� 
��     �a    �  �{ /B /Just L /Fields /Indent 0 /Text Paste (shortc    e-click the file to play it. ������    �   +�  �   in the Options, Preferences dialog, you can also doubl�  ust L /Fields /Indent 0 /Text Note: If you have specified�  ress F5, or click File, Play. ����u�  �  �� /P /J�  DVA. ����<"  O  �J /E /Just L /Fields /Indent 0 /Text P�   /Fields /Indent 0 /Text Open the file you wish to play in �   L /Fields /Indent 0 /Text OR������  Q  �L /E /Just L�  ht-click the file and click Play.��ql  .  �) /P /Just�   /Indent 0 /Text From a Windows Explorer window, simply rig�   11To play a file:���� 3  u  �p /B /Just L /Fields�   files.���� ˳  @  �; /4 /Just L /Fields /Indent 0 /Text�  lds /Indent 0 /Text ��DVA can play MVA files as well as DVA�  ent 0 /Text Playing a File�� �h  X  �S /P /Just L /Fie�   0 �� ��     � 9 �� �  8  �3 /1 /Just L /Fields /Ind�  lected text in the clipboard without deleting it. ����)��  ng through Windows is too slow or low in quality. ���� ��  .mva files to an MS-DOS Batch file. This is useful if playi�   L /Fields /Indent 0 /Text ��DVA can compile both .dva and �   /Indent 0 /Text Compiling a File�� ��  �  �� /P /Just�    � 0 �� ��     � 11 �� �  :  �5 /1 /Just L /Fields�  ling a File�� W�     �  �� 	g�     � Topic1�� 
��   �      �    �    �  ��A^     �  �� H~     � Compi�  Z  �m��E E  3 : O     � Topic@Compiling a File  ��  Y /Indent 0 /Width /Height�� �   �  �� /P /Just L /Field�  s /Indent 0 /Text Times New Roman12��The Edit menu�   (Alt+E) contains commands for working with text in the �  editing area. ���� �  z  �u /B /Just L /Fields /Indent �  0 /Text Cut (shortcut Ctrl+X) Deletes selected text and�   placed it in the clipboard. ���� �0  �  �{ /B /Just L /�  Fields /Indent 0 /Text Copy (shortcut Ctrl+C) Places sen�    D  �? /4 /Just L /Fields /Indent 0 /Text 11To compile       �   �J                                          �  le just by double-clicking it in Windows Explorer.��Q �  fied so in Options, Preferences, you can compile the fi�  P /Just L /Fields /Indent 0 /Text Note: If you have speci�  re you want to place the compiled file. �����A  �  �� /�  Just L /Fields /Indent 0 /Text Browse for the directory whe�  ss F6, or click File, Compile. ����\�  n  �i /E /�  A. ����#  R  �M /E /Just L /Fields /Indent 0 /Text Pre�  lds /Indent 0 /Text Open the file you wish to compile in DV�  ields /Indent 0 /Text OR������  T  �O /E /Just L /Fie�  to place the compiled file. ����&S  .  �) /P /Just L /F�  ds /Indent 0 /Text Browse for the directory where you want �  nd then click Compile. �����  n  �i /E /Just L /Fiel�  Text From a Windows Explorer window, right-click the file a�   a file: ���� �  y  �t /E /Just L /Fields /Indent 0 /n/  rap toggles word wrapping in the editing area. ������   Text New (shortcut Ctrl+N) clears the text area and let�  nd MVA files:�� ��  �  �� /B /Just L /Fields /Indent 0 /�  (Alt+F) contains the following items for working with DVA a�  s /Indent 0 /Text Times New Roman12��The File menu �  Y /Indent 0 /Width /Height�� �  �  �� /P /Just L /Field�  \FILEMENU.BMP /Macro /Play /Popup /Border 0 /Just L /Stack �  �� �y  �  �� /I /Jump /Link j:\HLP\WINHELP4\SOURCE\COMMON�  ��   3  �. /1 /Just L /Fields /Indent 0 /Text File Menu�  �� �y  �  �� /I /Jump /Link j:\HLP\WINHELP4\SOURCE\COMMON�  \VIEWMENU.BMP /Macro /Play /Popup /Border 0 /Just L /Stack �  Y /Indent 0 /Width /Height�� ��  ?  �: /P /Just L /Field�  s /Indent 0 /Text Times New Roman12���� �L  ~  �y /B�   /Just L /Fields /Indent 0 /Text Refresh (shortcut F5)    reloads the file list on the left hand side of the window.��  ��� ��  a  �\ /B /Just L /Fields /Indent 0 /Text Word W�  s you create a new file. You will be promted to save any ch  ve As... prompts you for a new filename for the open file.  e. ����49  i  �d /B /Just L /Fields /Indent 0 /Text Sa  If the file is untitled, you will be prompted for a filenam  Ctrl+S) saves the currently open file with its filename.    �  �� /B /Just L /Fields /Indent 0 /Text Save (shortcut   ayed later outside DVA or from DOS as you wish. ������   nt DVA or MVA file to an MS-DOS Batch file, which can be pl  Compile... (shortcut F7) allows you to export the curre	  tely. �����  �  �� /B /Just L /Fields /Indent 0 /Text 
  ay (shortcut F6) plays the currently opened file immedia  e. ����&+  n  �i /B /Just L /Fields /Indent 0 /Text Pl  l be promted to save any changes to the originally open fil  lets you open a previously written DVA or MVA file. You wil  st L /Fields /Indent 0 /Text Open... (shortcut Ctrl+O)   anges to the originally open file. ���� ��  �  �� /B /Ju    �����  �  �� /B /Just L /Fields /Indent 0 /Text Prin�  c  ����? �  0 7 L     � Topic@Saving a File  �  Y   � 0 �� ��   6  �1 /1 /Just L /Fields /Indent 0 /Text Op   P�     �  �� 	`�     �	 View Menu�� 
y�     � 0 �� �  ��   3  �. /1 /Just L /Fields /Indent 0 /Text View Menu   P�     �  �� 	`�     �	 Edit Menu�� 
y�     � 0 ��   ��   3  �. /1 /Just L /Fields /Indent 0 /Text Edit Menu  �� �y  �  �� /I /Jump /Link j:\HLP\WINHELP4\SOURCE\COMMON�  \EDITMENU.BMP /Macro /Play /Popup /Border 0 /Just L /Stack     changes. ������    � 13 ��a     �   ��      cut Alt+F4) closes DVA. You will be prompted to save any   B�  {  �v /B /Just L /Fields /Indent 0 /Text Exit (short  you to view and edit file properties in a dialog box����   /B /Just L /Fields /Indent 0 /Text Properties... allows   e specified in Options, Preferences.... �����X  u  �p  t (shortcut Ctrl+P) prints the file to the device or filn�   P�     �  �� 	`�     �	 File Menu�� 
y�     � 0 �� #  where the last string was found. Note that if you select F$  ind... again, any subsequent searches will take place from%   the beginning of the open file. ����GI  3 �./B /Just&   L /Fields /Indent 0 /Text Replace... (shortcut Ctrl+H)'   searches for all instances of a particular item of text an(  d replaces it with text you specify. If you select text wit�  hin the editing area before you select Replace, this text w�  with Inno-Setup, a freeware tool available from 1www.jrso)  GET� /Indent 0 /Text The setup program for DVA was created *  acroArg2 �Jump �HREF http:��www.jrsoftware.org �Anchor �TAR+  bX  �  �� /B /Just L /Fields 1�87�104��Macro �MacroArg1 �M,  reated with Windows Help Workshop version 4.03.0002.����4  s  o���9 �  . 5 J     � Topic@Search Menu  �          � 6 ��U�    �   ��                           enu�� S�     �  �� 	c�     � Options Menu�� 
�    "   (shortcut F3) re-executes the last find, beginning from     sion '.wad'. ����ĥ    � 6 ��<�    �   �� /  mp /Link j:\HLP\WINHELP4\SOURCE\COMMON\PROPDLG.BMP /Macro /5   �    �    �  ��<Y     �  �� Ct     � Search Men6  u�� R�     �  �� 	b�     � Search Menu�� 
}�     �7   0 �� ��   5  �0 /1 /Just L /Fields /Indent 0 /Text Searc8  h Menu�� ��  �  �� /I /Jump /Link j:\HLP\WINHELP4\SOURC9  E\COMMON\SEARCH~1.BMP /Macro /Play /Popup /Border 0 /Just L:   /Stack Y /Indent 0 /Width /Height�� �>  �  �� /P /Just ;  L /Fields /Indent 0 /Text Times New Roman12��The Sea<  rch menu (shortcut Alt+S) contains commands for finding =  and replacing text within the editing area: ���� ��  �  >  �� /B /Just L /Fields /Indent 0 /Text Find... (shortcut ?  Ctrl+F) displays a dialog box where you can search for a t@  ext string within the currently open DVA or MVA file. ����1   �   �/B /Just L /Fields /Indent 0 /Text Find Next2  n your sounds directory. DVA Wave Data files have the extenQ  Index (shortcut Shift+F1)displays the index page of the B  ile. ���� �  t  �o /B /Just L /Fields /Indent 0 /Text C   (shortcut F1) opens the contents page of the DVA help fD  �� �  s  �n /B /Just L /Fields /Indent 0 /Text ContentsE   (Alt+H) takes you to instant local and online help. ��F  s /Indent 0 /Text Times New Roman12��The Help menuG  Y /Indent 0 /Width /Height�� �  �  �� /P /Just L /FieldH  \HELPMENU.BMP /Macro /Play /Popup /Border 0 /Just L /Stack I  �� �y  �  �� /I /Jump /Link j:\HLP\WINHELP4\SOURCE\COMMONJ  ��   3  �. /1 /Just L /Fields /Indent 0 /Text Help MenuM  Menu Reference�� �!� T�1�File Menu�File Menu� �!� T�1�EdiN  t Menu�Edit Menu� �!� T�1�View Menu�View Menu� �!� T�1�SeO  arch Menu�Search Menu� �!�  T�1�Options Menu�Options Menu� �  �!� T�1�Help Menu�Help Menu� �!�# F�0�Keyboard Shortcut ReA  .wav), renaming it to a DVA Wave Data file and placing it i"`  DVA help file.�����  o  �j /B /Just L /Fields /Indent S  nt programs were created completely with freeware programs.T   Therefore, DVA is distributed for non-commercial use as frU  eeware, and it will remain that way. ���� �Y  R �M/B /V  Just L /Fields 1�138�161��Macro �MacroArg1 �MacroArg2 �JumpW   �HREF http:��www.basicguru.com�rapidq �Anchor �TARGET� /InX  dent 0 /Text The actual DVA program was written in Rapid-Q.Y   This is a freeware, object-oriented 32-bit compiler and inZ  terpreter. It is available from 1www.basicguru.com/rapidq[   and was created by William Yu.���� �  q  �l /B /Just \  L /Fields /Indent 0 /Text The CHM documentation was created]   with HTML Help Workshop version 4.74.����Y  y  �t /B -  /Just L /Fields /Indent 0 /Text The HLP documentation was c    �                                                       ^  information, etc. ������    � 7 ���    �   �_  0 /Text About... shows a dialog box containing copyright *R  Fields /Indent 0 /Text ��DVA and all its associated assistac    �    �    �  ��?\     �  �� Fz     � Compiled   Dialog�� U�     �  �� 	e�     � Compile Dialog�� 
�e  �     � 0 �� ��   8  �3 /1 /Just L /Fields /Indent 0 /Te�  xt Compile Dialog�� ��  �  �� /P /Just L /Fields /Inde    ol. See the Windows Help.�� ň    �    �        f  nt 0 /Text ��The file open dialog is a Windows common contrg  /Text Open Dialog�� �x  q  �l /P /Just L /Fields /Indeh   ��     � 3 �� ��   5  �0 /1 /Just L /Fields /Indent 0 i  g�� R�     �  �� 	b�     � Topic1�� 
}�     � 0 ��j   �    �    �  ��<Y     �  �� Ct     � Open Dialom  q  ���9 l  2 9 N     � Topic@Creation of DVA  � n     �    �    �  ��@]     �  �� G|     � Creatio  on of DVA�� V�     �  �� 	f�     � Topic1�� 
��    p   � 0 �� ��     � 7 �� �  9  �4 /1 /Just L /Fields /Ia  ndent 0 /Text Creation of DVA�� ��  �  �� /P /Just L /b  �  ����- �  1 8 M     � Topic@Compile Dialog  �      rtcut Reference� �                                         3  s /Indent 0 /Text Properties Dialog�� ��  �  �� /I /Jus      � 0 �� ��     � 4 �� �  ;  �6 /1 /Just L /Fieldt  erties Dialog�� X�     �  �� 	h�     � Topic1�� 
�� u  �    �    �    �  ��B_     �  �� I�     � Propv  �  ���0 �  4 ; P     � Topic@Properties Dialog  )   /Fields /Indent 0 /Text ��This dialog will prompt you whet    1 VHOBJECT22 VHOBJECT23 VHOBJECT24 VHOBJECT25 VHOBJECT26   D    �    �  ��7T     �  �� >w     � Save Changes Diz  alog�� M�     �  �� 	]�     � Topic1�� 
��     � 0    �� ��    � 3 �� ��    �    ��                |  ight information, acknowledgements and version information.}  xt Times New Roman12��The About dialog displays copyr~  out Dialog�� ��  �  �� /P /Just L /Fields /Indent 0 /Te   � 0 �� ��   6  �1 /1 /Just L /Fields /Indent 0 /Text Abnr  ference�� �!�> T�1�Keyboard Shortcut Reference�Keyboard Sho�  currently open file. ������  f  �a /B /Just L /Fields /�    O  �J /B /Just L /Fields /Indent 0 /Text F6: Plays the �  Indent 0 /Text Ctrl+O: Opens an existing file. ����SN�   Creates a new file. ������  L  �G /B /Just L /Fields /�  �� 6�  H  �C /B /Just L /Fields /Indent 0 /Text Ctrl+N:�  Arg2 /HREF /Anchor /TARGET /Fields /Text ��File Menu���  ink /Macro /Play /Popup /Just L /Indent 0 /MacroArg1 /Macro�   to access dialogs. ���� �J  �  �� /L /Jump File Menu /L�   ��These are all the keyboard shortcut commands you can use�  eference�� ԰  x  �s /P /Just L /Fields /Indent 0 /Text�   �@ /1 /Just L /Fields /Indent 0 /Text Keyboard Shortcut R�    � Topic1�� 
��     � 0 �� ��     � 26 �� �-  E �     � Keyboard Shortcut Reference�� b�     �  �� 	r�   �  erence  �    �    �    �  ��Li     �  �� S�   �  g  ����r &g  > E Z   &  �! Topic@Keyboard Shortcut Ref��  Indent 0 /Text F7: Displays a dialog to compile the curre�   ���� u  �  �{ /B /Just L /Fields /Indent 0 /Text Ctrl�   Places selected text on the clipboard without deleting it.�  ��f�  o  �j /B /Just L /Fields /Indent 0 /Text Ctrl+C:�  letes the selected text and places it on the clipboard. ���  �p  n  �i /B /Just L /Fields /Indent 0 /Text Ctrl+X: De�  2 /HREF /Anchor /TARGET /Fields /Text ��Edit Menu�����   /Macro /Play /Popup /Just L /Indent 0 /MacroArg1 /MacroArg�  to save changes. ����i�  �  �� /L /Jump Edit Menu /Link�  lds /Indent 0 /Text Alt+F4: Closes DVA. You are prompted �  ons | Set Print Output... �����]  b  �] /B /Just L /Fie�  P: Prints the file to the device or file specified in Opti�  ����W�  �  �� /B /Just L /Fields /Indent 0 /Text Ctrl+�  ile is untitled, you are prompted for a name and location. �  t 0 /Text Ctrl+S: Saves the currently open file. If the f�  ntly open file. �����`  �  �� /B /Just L /Fields /Inden�  +V: Inserts text on the clipboard into the editing area at�  ����	!�9  �  �� /B /Just L /Fields /Indent 0 /Text Ctrl+�   ;  �6 /B /Just L /Fields /Indent 0 /Text F3: Find Next. �  ialog allowing you to search for a text string. ���� >�
 �  /Just L /Fields /Indent 0 /Text Ctrl+F: Displays a Find d�  TARGET /Fields /Text ��Search Menu�����S
  u  �p /B �  pup /Just L /Indent 0 /MacroArg1 /MacroArg2 /HREF /Anchor /�  ��;�	  �  �� /L /Jump Search Menu /Link /Macro /Play /Po�  Text F5: Reloads file list on left hand side of window.���  View Menu�����5	  ^  �Y /B /Just L /Fields /Indent 0 /�  croArg1 /MacroArg2 /HREF /Anchor /TARGET /Fields /Text ���  p View Menu /Link /Macro /Play /Popup /Just L /Indent 0 /Ma�  ll text in the text editing area. ����~�  �  �� /L /Jum�    �Z /B /Just L /Fields /Indent 0 /Text Ctrl+A: Selects a�  /Indent 0 /Text Del: Deletes selected text. �����2  _�   the insertion point. ����y�  H  �C /B /Just L /Fields �  H: Displays Replace dialog so you can replace all instance�  le: These files are source files created by a program simi�  lar to DVA called MVA, and hence have the extension '.mva'.�   DVA has the ability to open, save, play and compile MVA fi�  les as you would a DVA file. MVA files are also plain ASCII�   text and can be edited with any text editor as well as fro�  m within DVA. ���� }�  V �Q/B /Just L /Fields /Indent �  0 /Text DVA Wave Data file: These are the sound bites whi�  ch are put together to make an announcement. You can add yoP  ur own simply by creating an uncompressed wave-sound file (    +F1: Displays Help index.��%�^    �   &'W       �  ����
$BN  H  �C /B /Just L /Fields /Indent 0 /Text Shift�  s /Indent 0 /Text F1: Displays Help contents and topics. �  ds /Text ��Help Menu����
#��  S  �N /B /Just L /Field�   /L /Jump /Link /Macro /Play /Popup /Just L /Indent 0 /Fiel�  s of particular text with different text. ����	"\�  Y  �T"�  3  m �h/B /Just L /Fields /Indent 0 /Text MVA Source fi�   �    �    �  ��<Y     �  �� Cw     � Save As Di�  �  ����- �  . 5 J     � Topic@Save Dialog  �   k  �   ���- �  . 5 J     � Topic@Open Dialog  �   �  �  <���6 �  - 4 I     � Topic@File Types  �    �  �    �    �  ��;X     �  �� Br     �
 File Types�  �� Q�     �  �� 	a�     �
 File Types�� 
{�     � 0 �  �� ��   4  �/ /1 /Just L /Fields /Indent 0 /Text File Typ�  es�� �t  }  �x /P /Just L /Fields /Indent 0 /Text Time�  s New Roman12��DVA has several related file types. The�  y are listed here. ���� ��  < �7/B /Just L /Fields /In�  dent 0 /Text DVA Source file: These files are what you cr�  eate when you write a source and then save it. They have th�  e extension '.dva'. These files are ASCII text so you can u�  se any non-formatting text editor such as Windows Notepad t�  o edit them, besides editing them from within DVA. ���� �"�  alog�� R�     �  �� 	b�     � Save Dialog�� 
��    �  �  ���3 �  / 6 K     � Topic@Options Menu  �  K   P�     �  �� 	`�     �	 Help Menu�� 
y�     � 0 �� �      �    �  ��:W     �  �� Ap     �	 Help Menu���  �  �J��9 �  , 3 H     � Topic@Help Menu  �    �     3 �� ��    �    ��                              E  eating a new file, if the current file has been modified si�  nce the last save. Click Yes to save changes, No to rejY  anges�� ��  �  �� /I /Jump /Link j:\HLP\WINHELP4\SOURCE        � 3 �� �    �   ��                        �   is a Windows common control. See the Windows help.�� £�  nt 0 /Text Times New Roman12��The file compile dialog�  Windows common control. See the Windows help.�� ��    ��  Text Times New Roman12��The file save-as dialog is a �  ve As Dialog�� ��  �  �� /P /Just L /Fields /Indent 0 /�   � 0 �� ��   8  �3 /1 /Just L /Fields /Indent 0 /Text Sa0    �    �    �  ��=Z     �  �� Dv     � Options M�  Indent 0 /Text Version History�� �I  5 �0/P /Just L �   � 0 �� ��     � 14 �� �	  9  �4 /1 /Just L /Fields /�  n History�� V�     �  �� 	f�     � Topic1�� 
��    �     �    �    �  ��@]     �  �� G|     � Versio�  �  r7��N t  2 9 N     � Topic@Version History  �     !�  !�  !�  !�  !�  !�                                     !      �    �  ��:W     �  �� Ap     �	 File Menu���  	  B���K �  , 3 H     � Topic@File Menu  �    �    rea. ����ı    � 9 ��-�    �   ��               �    �  ��:W     �  �� Ap     �	 View Menu���  �   ���6 �  , 3 H     � Topic@View Menu  �    �      �    �  ��:W     �  �� Ap     �	 Edit Menu���  �  (���? �  , 3 H     � Topic@Edit Menu  �    ��  ill automatically be entered into the Replace edit box. ��    ��Z    � 7 ��j    �   Rc                 n   /Fields /Indent 0 /Text ��v4.00��Fourth generation. Opera   new one-click DVA Autoplay and Upgrade! Now you can upgrad�  imation with sound too! Now for the most inportant upgrade,�  e DVA example files. Included a brand new logo and title an�   More sounds from Sydney, as well as Brisbane now. Even mor�  sn't have to be searched through and edited by the program.�  eds up the upgrade process, as the entire wads.dat file doe�  tomised data is stored in the file user.dat, which also spe�  xt v3.0x��Even greater user customisability. The user-cus�   4 above.���� $  M �H/P /Just L /Fields /Indent 0 /Te�   Fourth generation beta��Fourth generation beta for version�  � ��  x  �s /P /Just L /Fields /Indent 0 /Text v0.40b -�  ck and ability to compile MVA/DVA files to BATch files.����  ck-builder, customisable shell integration, enhanced playba�  index files. Extensive MVA support, built in editor and qui�  tes fully in Windows 32-bit GUI. No more DOS! Also no more n  e or play DVA files from anywhere. Right-click context menu   DVA data (.wad), and a fancy new icon for it! Worked out h  ludes more station data. Created a unique file type for the  o have found a setup program THAT ACTUALLY WORKS!! Also inc  �&/P /Just L /Fields /Indent 0 /Text v2.03��Now I seem t   and to let the user add his/her own sounds.������  +   the net. Created a new play engine, to make upgrades easier   run-time compiler, after recovering a corrupted file from    startup. Also added some more DVA example files. Abolished	  ent 0 /Text v2.10��Included a splash screen to display at
  ed icons.dll file.����-�  6 �1/P /Just L /Fields /Ind  ields /Indent 0 /Text v2.11��Added more sounds, and updat   Explorer Shell integration.�����J  a  �\ /P /Just L /F   beta for third generation (3.x) version, implementing full  dent 0 /Text v0.30b - Third generation beta��Experimental   in Explorer added.����R�  �  �� /P /Just L /Fields /In�   ow to use setup compression, reducing the file size by 40%.!  l data yet though.����	��  l  �g /P /Just L /Fields /Ind  n experimental. Brightened up the interface. Don't have ful  /Just L /Fields /Indent 0 /Text v0.20 - Second beta��Agai  n uninstall, and an internet shortcut.����Z  �  �� /P   hap during downloading. Also added some snazzy new icons, a  file, and broke up the volumes into pieces in case of a mis   source files. Added a Setup executable to replace the zip   ugs in recognising 'Wentworth Falls' and 'Milsons Point' in  ext v2.00 - First full release��No full data, but fixed b   zip file.�����p  s �n/P /Just L /Fields /Indent 0 /T   setup creator, the method of distribution is reverted to a  lds /Indent 0 /Text v2.01��Due to serious faults with the  ams, and was not released.������	  �  �� /P /Just L /Fie  ��Version created, but even more problems with setup progr  ����SQ	  �  �� /P /Just L /Fields /Indent 0 /Text v2.020  ent 0 /Text v0.10 - First beta��Experimental version. Min1   ��     � 5 �� ��   5  �0 /1 /Just L /Fields /Indent 0 "  g�� R�     �  �� 	b�     � Topic1�� 
}�     � 0 ��#   �    �    �  ��<Y     �  �� Ct     � Find Dialo$  �  b���3 �  . 5 J     � Topic@Find Dialog  �   4    �    �    �  ��?\     �  �� Fz     � Replace&  0  ���0 �  1 8 M     � Topic@Replace Dialog  �  �  \COMMON\SAVECH~1.BMP /Macro /Play /Popup /Border 0 /Just L (  /Stack Y /Indent 0 /Width /Height�� ��   �/P /Just L    ved as a DVA file.�� �    �   ��               *   properties cannot be added or changed until the file is sa+  on about the file. If the file being edited is an MVA file,,  e file properties dialog allows you edit and view informati-  ight�� ј  �  �� /P /Just L /Fields /Indent 0 /Text ��Th.  Play /Popup /Border 0 /Just L /Stack Y /Indent 0 /Width /He    imal data included.����	y�    �   �            @  /Text Find Dialog�� ��  �  �� /I /Jump /Link j:\HLP\WIA  ent 0 /Text Replace Dialog�� ��  �  �� /I /Jump /Link 2   0 �� ��     � 4 �� �  8  �3 /1 /Just L /Fields /Ind3   Dialog�� U�     �  �� 	e�     � Topic1�� 
��     �    �                                                      5  st L /Stack Y /Indent 0 /Width /Height����    �   6  4\SOURCE\COMMON\NFDLG.BMP /Macro /Play /Popup /Border 0 /Ju7  ing are found.�� �  �  �~ /I /Jump /Link j:\HLP\WINHELP8  ialog will be shown when no more occurences of the text str9  nu to find further occurences of the text string.����This d:  will be highlighted. Click Find Next from the Search me;  the string and click Find to search. The first occurence <  ws you to search the current file for a text string. Enter =  n/P /Just L /Fields /Indent 0 /Text ��The Find dialog allo>  r 0 /Just L /Stack Y /Indent 0 /Width /Height�� �
  s �?  NHELP4\SOURCE\COMMON\FINDDLG.BMP /Macro /Play /Popup /Borde"P  j:\HLP\WINHELP4\SOURCE\COMMON\REPLAC~1.BMP /Macro /Play /PoQ      �    �  ��:W     �  �� Ap     �	 Locations��B  B  1>��0 �  , 3 H     � Topic@Locations  �    �s  �  ���0 �  ) 0 E     � Topic@Topic1  �    �  x  her to save changes when closing DVA, opening a file, or crG  �  ���- �  / 6 K     � Topic@About Dialog  �  H    �    �    �  ��=Z     �  �� Dv     � About Dia�  log�� S�     �  �� 	c�     � About Dialog�� 
�        ly be placed in the dialog.�� '    �   �       I   area before selecting Replace, the text will automaticalJ   with, and click OK. If you highlight text in the editingK  replace and the string you want to replace the first stringL  ng with another text  string. Enter the string you want to M  e dialog allows you to replace all instances of a text striN  �  v �q/P /Just L /Fields /Indent 0 /Text ��The ReplacO  pup /Border 0 /Just L /Stack Y /Indent 0 /Width /Height�� "`   P�     �  �� 	`�     � Topic1�� 
y�     � 0 �� ��a  0 /Just L /Stack Y /Indent 0 /Width /Height�� �d  �  �� R  LP4\SOURCE\COMMON\APPEAR~1.BMP /Macro /Play /Popup /Border S  ext Appearance�� ��  �  �� /I /Jump /Link j:\HLP\WINHET  ��     � 4 �� ��   4  �/ /1 /Just L /Fields /Indent 0 /TU  �� Q�     �  �� 	a�     � Topic1�� 
{�     � 0 �� V  �    �    �  ��;X     �  �� Br     �
 AppearanceW  }  �f��0 �  - 4 I     � Topic@Appearance  �    {   �� ��   6  �1 /1 /Just L /Fields /Indent 0 /Text Save Ch    urces and printer output.�� �9    �    �2        Z  ws you to set and view the default locations for sounds, so[  /Just L /Fields /Indent 0 /Text ��The Locations dialog allo\  Just L /Stack Y /Indent 0 /Width /Height�� �)  �  �� /P ]  \SOURCE\COMMON\LOCATI~1.BMP /Macro /Play /Popup /Border 0 /^  t Locations�� ��  �  �� /I /Jump /Link j:\HLP\WINHELP4_       � 4 �� ��   3  �. /1 /Just L /Fields /Indent 0 /Texp  /P /Just L /Fields /Indent 0 /Text ��In the Appearance sect�  ect changes since the last save.�� ��    � 4 �� ��        �    �I                                            c   MVA file is double-clicked in Windows Explorer.�� �P  d  es dialog, you can specify the default action when a DVA ore  lds /Indent 0 /Text ��In the Shell section of the Preferencf  k Y /Indent 0 /Width /Height�� �@  �  �� /P /Just L /Fieg  ON\SHELLDLG.BMP /Macro /Play /Popup /Border 0 /Just L /Stach  �� �{  �  �� /I /Jump /Link j:\HLP\WINHELP4\SOURCE\COMMi   4 �� ��   /  �* /1 /Just L /Fields /Indent 0 /Text Shellj    �  �� 	\�     � Topic1�� 
q�     � 0 �� ��     �k    �    �  ��6S     �  �� =h   
  � Shell�� Lx   l  Y  ����0 �  ( / D     � Topic@Shell  �    �       font used in the editor.�� t    �   �m        n  relating to how DVA looks including toolbar options and theo  ion of the Preferences dialog, you can set various options ob    �   ��                                                                                                          r                                                                 ve.�� �    �   ��                              t   to save changes, No to reject changes since the last sau  rent file has been modified since the last save. Click Yesv  ing DVA, opening a file, or creating a new file, if the curw  is dialog will prompt you whether to save changes when closx  ight�� ��   �/P /Just L /Fields /Indent 0 /Text ��Thy  Play /Popup /Border 0 /Just L /Stack Y /Indent 0 /Width /Hez  p /Link j:\HLP\WINHELP4\SOURCE\COMMON\SAVECH~1.BMP /Macro /{  ields /Indent 0 /Text Save Changes�� Ğ  �  �� /I /Jum|  
��     � 0 �� ��     � 4 �� �  6  �1 /1 /Just L /F}  ve Changes Dialog�� Z�     �  �� 	j�     � Topic1�� ~    �    �    �    �  ��Da     �  �� K�     � Sa  �  _��0 �  6 = R     � Topic@Save Changes Dialog