���Z     @     IH        <&                                                                                                !   �   zY 	   ,          � Project@Options� -�   !�     7   |+ 	   -          � File@@Version2.1  � 1.2 =   @                                                          1   �   TOPIC VERSION OBJARRAY BROWSE_SEQUENCE BUILD_TAG CONTEX    link viewHandles 7                                            _ISECT_iterator _AE_Sorter _AE_mark _SysInfoFlags _outside_   Metafile VbPicture VbVarArray VeRec ViewEngine WinImage _AE   r VB_Historian VB_View VbCurrency VbDibBitmap VbFixArray Vb	   ng SystemDatabase TextFileDatabase TrashCollector TreeWalke
   Real RecordMark RuleSpecifier SchemaEngine SmartString Stri   adStream NamedData NamedMonad NilMonad Number Presentation    Dictionary Integer LogStream Monad MonadArray MonadFile Mon   tion Bcd36 Boolean ClassDesc ClassMethod ComboElement Date    Set AdRec AeAccessSet AgilityDatabase ArrayDatabase Associa   ]  YAccessCombo AccessEngine AccessItem AccessRule AccessH	 Z                   .       *       (       %       ]             \                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �0    !� BuildAll!� 0!� License Agreement!�$ Copyright � 1999#   , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 ,x     20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12    "", , , , (192,192,192), 0!�- "", ( 64, 64, 832, 832), , $   i  �� 	   -          � F1ProjectWindows:-�   !�    �  !�  !�  !�  !�  !�  !�  !�                              &     !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !�  !'   �   �4 	   -          � F1ProjectButtonsb -�   !�    �                                                          )   :   �� 	   .          � F1ProjectGlossary
 -�   !     !�  !�  !�  !�  !�  !�                                    +   bin\imagemap\!� d:\DVADev\hlp\!� _!�  !�  !�  !�  !�  !� ,    !� common!� 0!� 0!� 1!� 1!� 0!�  www.domain.com\cgi--   �   n	 	   0          � Project@OptionsHTML� -�      No!�  !� License Agreement!� 1!�  0!�  !�  !�           /   -2001 Jonathan Boles!�  !�  !�  !� 0!�  !�  !� 0!� 0!� B>   T_STRING HELP_MACRO KEYWORDS TOPIC_TITLE NOTE FILENAME PAGE3   , !�G Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 ,4    -1 ,  0 , None , !�G Heading , Arial ,  14 ,  120 ,  90 , 5    60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  146    ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Headi7   ng , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , 8   None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 ,  9   20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 , :    120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub Head;   ing , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 ,<    None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 , ?    20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12 ,                                                                   WIDTH VHOBJECT0 VHOBJECT1 VHOBJECT2 VHOBJECT3              @     120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub Hea"   ding , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 
2   Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None C   l ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�D   F Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,E     0 , None , !�E Title , Arial ,  18 ,  120 ,  90 ,  60 ,  F   20 ,  0 , -1 ,  0 , None , !�E Title , Arial ,  18 ,  120 ,G     90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�E Title , Arial H   ,  18 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�E I   Title , Arial ,  18 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0J    , None , !�E Title , Arial ,  18 ,  120 ,  90 ,  60 ,  20 K   ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14 ,  120 , L    90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , ArialM    ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�GN    Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,O     0 , None , !�G Heading , Arial ,  14 ,  120 ,  90 ,  60 ,P     20 ,  0 , -1 ,  0 , None , !�G Heading , Arial ,  14 ,  1A   20 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�G Heading , NB   ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�F Normal , Ariaa    a different license agreement signed by the author your usR    and conditions before using this software. Unless you haveS   mission.������You should carefully read the following termsT   ethell, Paul McCabe and Winston Yang.��Sounds used with perU   999 - 2001 Jonathan Boles��Sounds copyright Glenn Jackson-BV   Fields /Indent 0 /Text Times New Roman12��Copyright 1W   ent 0 /Text License Agreement�� �F  3 �./P /Just L /X   ent�� 
��     � 0 �� �  ;  �6 /1 /Just L /Fields /IndY   nse Agreement�� X�     �  �� 	h�     � License AgreemZ   �    �    �    �  ��B_     �  �� I�     � Lice[   p  -��-   4 ; P     � Topic@License Agreement  ^   �)  �� 	   ,          � F1ProjectStyle2�)-�  � !�F_    Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 , `    0 , None , !�F Normal , Arial ,  10 ,  120 ,  90 ,  20 ,  Q   20 ,  0 ,  0 ,  0 , None , !�F Normal , Arial ,  10 ,  120 �p   e of this software indicates your acceptance of this licensq   ISTRIBUTION ����You are not licensed to make copies of theb   not reverse, disassemble, decompiler, or alter DVA.������Dc   he DVA software is strictly not to be distributed. You may d   s you wish. DVA files may be distributed as you like, but te   low, you are licensed to use this software without charge af   ���USE ����This is free software. Subject to the terms beg   thor will be limited exclusively to product replacement.���h    entire risk of using the software, any liability of the aui   anties whether expressed or implied. ��The user assumes thej   ties as to performance or merchantability or any other warrk   files are supplied on an "as is" basis. There are no warranl   LAIMER OF WARRANTY ����This software and the accompanying m   accept this license agreement, click Cancel now.������DISCn    version or release of DVA. ��If you do not agree with and o   e agreement and warranty. This license agreement covers anyv�    DVA software and documentation except as stated below.��Yo�   0 , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60r   eading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  s    ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub Ht   ,  20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  12u    , None , !�K Sub Heading , Arial ,  12 ,  120 ,  90 ,  60 v   ading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0w   ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub He  This agreement shall be governed by laws of Australia.����y   e original Setup executable file.������GOVERNING LAW ����z   up purposes. Even then it is preferred if this backup is th{    software, including .wad files is allowed, solely for back|   Bethell, Paul McCabe and Winston Yang.��ONE copy of the DVA}   h DVA. Copyright of these files remains with Glenn Jackson-~   breaching copyright on ANY .wad files that are included wit   u are VERY STRICTLY prohibited from copying or otherwise ��    ,  20 ,  0 , -1 ,  0 , None , !�K Sub Heading , Arial ,  1�   0 ,  0 ,  0 , None , !�O Image Paragraph , Arial ,  10 ,  1�    Image Paragraph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  �    ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�O�   0 ,  20 ,  0 ,  0 ,  0 , None , !�O Image Paragraph , Arial�    None , !�O Image Paragraph , Arial ,  10 ,  120 ,  90 ,  2�   aph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 ,�    ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�O Image Paragr�    ,  0 ,  0 ,  0 , None , !�I Paragraph , Arial ,  10 ,  120�   None , !�I Paragraph , Arial ,  10 ,  120 ,  90 ,  20 ,  20�   ph , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , �     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�I Paragra�   ,  20 ,  0 ,  0 ,  0 , None , !�I Paragraph , Arial ,  10 ,�    0 , None , !�I Paragraph , Arial ,  10 ,  120 ,  90 ,  20 �   Heading , Arial ,  12 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 , �   2 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�K Sub ��   20 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnote ,�   0 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Numb�   ,  0 ,  0 ,  0 , None , !�R Numbered List Item , Arial ,  1�    Bulleted List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 �    ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R�     20 ,  0 ,  0 ,  0 , None , !�R Bulleted List Item , Arial�   , !�R Bulleted List Item , Arial ,  10 ,  480 ,  90 ,  20 ,�   Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None �    20 ,  20 ,  0 ,  0 ,  0 , None , !�R Bulleted List Item , �   None , !�R Bulleted List Item , Arial ,  10 ,  480 ,  90 , �   ote , Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , �    ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footn�    20 ,  20 ,  0 ,  0 ,  0 , None , !�G Footnote , Arial ,  8�     0 ,  0 , None , !�G Footnote , Arial ,  8 ,  120 ,  90 , �   , !�G Footnote , Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,�    Arial ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None ��   ered List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 �   10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�K Im�   0 ,  20 ,  10 ,  0 ,  0 , None , !�K Image Link , Arial ,  �     0 , None , !�K Image Link , Arial ,  10 ,  120 ,  90 ,  2�   ge Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,�   0 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�K Ima�    ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�E Link , Arial ,  1�     10 ,  0 ,  0 , None , !�E Link , Arial ,  10 ,  120 ,  90�    , None , !�E Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,�   Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0�     10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 ,  0 , None , !�E �     90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Link , Arial ,�   ,  0 , None , !�R Numbered List Item , Arial ,  10 ,  480 ,�   List Item , Arial ,  10 ,  480 ,  90 ,  20 ,  20 ,  0 ,  0 �   480 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Numbered �   ,  0 ,  0 , None , !�R Numbered List Item , Arial ,  10 ,  �   age Link , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  10 ,  0 �    ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Glossary Term , Ar�    ,  0 , None , !�M Index Heading , Arial ,  14 ,  120 ,  90�   ex Heading , Arial ,  14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1�   14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Ind�   ,  20 ,  0 , -1 ,  0 , None , !�M Index Heading , Arial ,  �    None , !�M Index Heading , Arial ,  14 ,  120 ,  90 ,  20 �   ing , Arial ,  14 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 ,�   20 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�M Index Head�    ,  20 ,  0 ,  0 ,  0 , None , !�E Index , Arial ,  10 ,  1�    0 ,  0 , None , !�E Index , Arial ,  10 ,  120 ,  90 ,  20�    , !�E Index , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �    Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None�     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Index ,�   20 ,  20 ,  10 ,  0 ,  0 , None , !�E Index , Arial ,  10 ,�   ,  0 , None , !�K Image Link , Arial ,  10 ,  120 ,  90 ,  J�   ial ,  12 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , �   -1 ,  0 , None , !�P Glossary Heading , Arial ,  14 ,  120 �   sary Heading , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , �   0 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�P Glos�     0 ,  0 ,  0 , None , !�S Glossary Definition , Arial ,  1�   lossary Definition , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,�     10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�S G�   0 ,  0 ,  0 ,  0 , None , !�S Glossary Definition , Arial ,�   S Glossary Definition , Arial ,  10 ,  120 ,  90 ,  20 ,  2�   l ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !��     20 ,  0 , -1 ,  0 , None , !�S Glossary Definition , Aria�   None , !�M Glossary Term , Arial ,  12 ,  120 ,  90 ,  20 ,�   rm , Arial ,  12 ,  120 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , �   0 ,  90 ,  20 ,  20 ,  0 , -1 ,  0 , None , !�M Glossary Te�    0 , -1 ,  0 , None , !�M Glossary Term , Arial ,  12 ,  12�   !�M Glossary Term , Arial ,  12 ,  120 ,  90 ,  20 ,  20 , N�   ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�P Glossary Head�     120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�E Table ,�    20 ,  20 ,  0 ,  0 ,  0 , None , !�E Table , Arial ,  10 ,�    ,  0 ,  0 , None , !�E Table , Arial ,  10 ,  120 ,  90 , �   one , !�E Table , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0�   urier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  5 ,  0 ,  0 , N�    90 ,  20 ,  20 ,  5 ,  0 ,  0 , None , !�P Button Bar , Co�    ,  0 , None , !�P Button Bar , Courier New ,  10 ,  120 , �    Bar , Courier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  5 ,  0�   ,  120 ,  90 ,  20 ,  20 ,  5 ,  0 ,  0 , None , !�P Button�   ,  5 ,  0 ,  0 , None , !�P Button Bar , Courier New ,  10 �   �P Button Bar , Courier New ,  10 ,  120 ,  90 ,  20 ,  20 �   al ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 , None , !�   60 ,  20 ,  0 , -1 ,  0 , None , !�P Glossary Heading , Ari�    None , !�P Glossary Heading , Arial ,  14 ,  120 ,  90 ,  �   ing , Arial ,  14 ,  120 ,  90 ,  60 ,  20 ,  0 , -1 ,  0 ,
�    Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None�    ,  440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�D Line �     10 ,  0 ,  0 ,  0 , None , !�L Outline Leaf , Arial ,  10�    None , !�L Outline Leaf , Arial ,  10 ,  440 ,  90 ,  10 ,�   eaf , Arial ,  10 ,  440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 ,�   440 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline L�    ,  0 ,  0 ,  0 , None , !�L Outline Leaf , Arial ,  10 ,  �   e , !�L Outline Leaf , Arial ,  10 ,  440 ,  90 ,  10 ,  10�   , Arial ,  10 ,  120 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , Non�   ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline Node �   0 ,  0 ,  0 , None , !�L Outline Node , Arial ,  10 ,  120 �   !�L Outline Node , Arial ,  10 ,  120 ,  90 ,  10 ,  10 ,  �   ial ,  10 ,  120 ,  90 ,  10 ,  10 ,  0 ,  0 ,  0 , None , �   0 ,  10 ,  10 ,  0 ,  0 ,  0 , None , !�L Outline Node , Ar�    0 ,  0 , None , !�L Outline Node , Arial ,  10 ,  120 ,  9�    , !�E Table , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , B   , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , Non  m Object , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20 ,  0�    8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R For�    ,  0 ,  0 ,  0 , None , !�R Form Object , MS Sans Serif , �   R Form Object , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20�   ial ,  10 ,  120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !��    120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 , None , !�C Image , Ar�     0 ,  0 ,  0 ,  0 ,  0 , None , !�C Image , Arial ,  10 , �   0 ,  0 ,  0 , None , !�C Image , Arial ,  10 ,  120 ,  90 ,�   , None , !�C Image , Arial ,  10 ,  120 ,  90 ,  0 ,  0 ,  �    Image , Arial ,  10 ,  120 ,  90 ,  0 ,  0 ,  0 ,  0 ,  0 �    ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�C�    ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�D Line , Arial�   ,  20 ,  0 ,  0 ,  0 , None , !�D Line , Arial ,  10 ,  120�    0 ,  0 , None , !�D Line , Arial ,  10 ,  120 ,  90 ,  20 �   e , !�D Line , Arial ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 , �   ,  0 ,  0 , None , !�R Form Object , MS Sans Serif ,  8 ,   4 "Glossary", ( 0, 0, 511, 1023), , , (192,192,192), 0!�3 "  192), 0!�. "", ( 0, 511, 1023, 511), , , (192,192,192), 0!�  , (192,192,192), 0!�, "", ( 0, 0, 1023, 511), , , (192,192,     !�  !�* T�0�License Agreement�License Agreement� �         k   �l 	   1          � F1ProjectContentList8 -�      20 ,  0 ,  0 ,  0 , None , !�                                 !�Q Mono Spaced , Courier New ,  10 ,  120 ,  90 ,  20 ,     New ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None ,	   20 ,  20 ,  0 ,  0 ,  0 , None , !�Q Mono Spaced , Courier
   None , !�Q Mono Spaced , Courier New ,  10 ,  120 ,  90 ,   Courier New ,  10 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 ,    90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�Q Mono Spaced ,    ,  0 , None , !�Q Mono Spaced , Courier New ,  10 ,  120 ,  ect , MS Sans Serif ,  8 ,  120 ,  90 ,  20 ,  20 ,  0 ,  0   120 ,  90 ,  20 ,  20 ,  0 ,  0 ,  0 , None , !�R Form Obj   Index", ( 511, 0, 511, 1023), , , (192,192,192), 0!�  !�  !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �W    � 3 �� g    �   O`                       �  !�  !�                                                  